module main

import erlang

fn main() {
	erlang.main()
}
